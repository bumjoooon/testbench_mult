module(mult_if _if);

assign _if.y = _if.a * _if.b;

endmodule
